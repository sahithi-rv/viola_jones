package IFC; 

// Multiplier IFC

import constants::*;

interface VJ_ifc;
    method Action  start (Bool x);
    method Pixels  result();
    
endinterface
        
endpackage